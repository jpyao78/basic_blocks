module clk_mux(
input i_clk0,
input i_clk1,
input i_sel,//0:o_clk= i_clk0;1:o_clk=i_clk1
output o_clk
);



endmodule
